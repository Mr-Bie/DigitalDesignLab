module dec4_16 (x,en,y);
input [0:3]x;
input en;
output reg [15:0]y;
always @(x,en)
case(x)
	4'b0000: y = 16'b1111111111111110;
	4'b0001: y = 16'b1111111111111101;
	4'b0010: y = 16'b1111111111111011;
	4'b0011: y = 16'b1111111111110111;
	4'b0100: y = 16'b1111111111101111;
	4'b0101: y = 16'b1111111111011111;
	4'b0110: y = 16'b1111111110111111;
	4'b0111: y = 16'b1111111101111111;
	4'b1000: y = 16'b1111111011111111;
	4'b1001: y = 16'b1111110111111111;
	4'b1010: y = 16'b1111101111111111;
	4'b1011: y = 16'b1111011111111111;
	4'b1100: y = 16'b1110111111111111;
	4'b1101: y = 16'b1101111111111111;
	4'b1110: y = 16'b1011111111111111;
	default: y = 16'b0111111111111111;
endcase
endmodule

